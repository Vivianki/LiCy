-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition"
-- CREATED		"Sat Sep 24 23:51:51 2016"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY RSencoder IS 
	PORT
	(
		Clock :  IN  STD_LOGIC;
		count :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		Output :  OUT  STD_LOGIC_VECTOR(0 TO 3);
		reg1 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		reg2 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		reg3 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		reg4 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		saida_AND :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		saidaMul :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END RSencoder;

ARCHITECTURE bdf_type OF RSencoder IS 

COMPONENT sinalcontrole
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 control : OUT STD_LOGIC;
		 count : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT scale_clock_100khz
	PORT(clk_50Mhz : IN STD_LOGIC;
		 rst : IN STD_LOGIC;
		 clk_100kHz : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT gf_mult
	PORT(x : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 y : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register4b
	PORT(ld : IN STD_LOGIC;
		 clr : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 d : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT gf_sum
	PORT(a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 b : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 c : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT and4x1
	PORT(b : IN STD_LOGIC;
		 a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 c : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux2x1
GENERIC (NB : INTEGER
			);
	PORT(Sel : IN STD_LOGIC;
		 I0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 I1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 O : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT static_13
	PORT(		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT static_4
	PORT(		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT static_14
	PORT(		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT static_8
	PORT(		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT static_1
	PORT(		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT static_0
	PORT(		 o : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC_VECTOR(3 DOWNTO 0);


BEGIN 
reg1 <= SYNTHESIZED_WIRE_55;
reg2 <= SYNTHESIZED_WIRE_63;
reg3 <= SYNTHESIZED_WIRE_65;
reg4 <= SYNTHESIZED_WIRE_77;
saida_AND <= SYNTHESIZED_WIRE_74;
saidaMul <= SYNTHESIZED_WIRE_14;
SYNTHESIZED_WIRE_73 <= '0';
SYNTHESIZED_WIRE_75 <= '1';
SYNTHESIZED_WIRE_78 <= "1111";



b2v_inst : sinalcontrole
PORT MAP(clk => SYNTHESIZED_WIRE_72,
		 reset => SYNTHESIZED_WIRE_73,
		 control => SYNTHESIZED_WIRE_76,
		 count => count);


b2v_inst1 : scale_clock_100khz
PORT MAP(clk_50Mhz => Clock,
		 rst => SYNTHESIZED_WIRE_73,
		 clk_100kHz => SYNTHESIZED_WIRE_72);


b2v_inst10 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_4,
		 o => SYNTHESIZED_WIRE_62);


b2v_inst11 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_6,
		 o => SYNTHESIZED_WIRE_14);


b2v_inst12 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_10,
		 q => SYNTHESIZED_WIRE_24);


b2v_inst13 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_14,
		 q => SYNTHESIZED_WIRE_55);


b2v_inst14 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_18,
		 q => SYNTHESIZED_WIRE_63);


b2v_inst15 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_22,
		 q => SYNTHESIZED_WIRE_65);



b2v_inst19 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_23,
		 b => SYNTHESIZED_WIRE_24,
		 c => SYNTHESIZED_WIRE_37);


b2v_inst2 : and4x1
PORT MAP(b => SYNTHESIZED_WIRE_76,
		 a => SYNTHESIZED_WIRE_26,
		 c => SYNTHESIZED_WIRE_74);


b2v_inst20 : mux2x1
GENERIC MAP(NB => 4
			)
PORT MAP(Sel => SYNTHESIZED_WIRE_76,
		 I0 => SYNTHESIZED_WIRE_77,
		 I1 => SYNTHESIZED_WIRE_78,
		 O => Output);


b2v_inst21 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_30,
		 b => SYNTHESIZED_WIRE_31,
		 c => SYNTHESIZED_WIRE_41);


b2v_inst22 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_32,
		 b => SYNTHESIZED_WIRE_33,
		 c => SYNTHESIZED_WIRE_45);



b2v_inst24 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_37,
		 q => SYNTHESIZED_WIRE_31);


b2v_inst25 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_41,
		 q => SYNTHESIZED_WIRE_33);


b2v_inst26 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_45,
		 q => SYNTHESIZED_WIRE_47);


b2v_inst27 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_46,
		 b => SYNTHESIZED_WIRE_47,
		 c => SYNTHESIZED_WIRE_51);


b2v_inst28 : register4b
PORT MAP(ld => SYNTHESIZED_WIRE_75,
		 clr => SYNTHESIZED_WIRE_73,
		 clk => SYNTHESIZED_WIRE_72,
		 d => SYNTHESIZED_WIRE_51,
		 q => SYNTHESIZED_WIRE_77);


b2v_inst29 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_53,
		 o => SYNTHESIZED_WIRE_23);


b2v_inst3 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_54,
		 b => SYNTHESIZED_WIRE_55,
		 c => SYNTHESIZED_WIRE_18);


b2v_inst30 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_57,
		 o => SYNTHESIZED_WIRE_30);


b2v_inst31 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_59,
		 o => SYNTHESIZED_WIRE_32);


b2v_inst32 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_61,
		 o => SYNTHESIZED_WIRE_46);


b2v_inst33 : static_13
PORT MAP(		 o => SYNTHESIZED_WIRE_6);


b2v_inst34 : static_13
PORT MAP(		 o => SYNTHESIZED_WIRE_53);


b2v_inst35 : static_13
PORT MAP(		 o => SYNTHESIZED_WIRE_61);


b2v_inst36 : static_4
PORT MAP(		 o => SYNTHESIZED_WIRE_71);


b2v_inst37 : static_14
PORT MAP(		 o => SYNTHESIZED_WIRE_4);


b2v_inst38 : static_8
PORT MAP(		 o => SYNTHESIZED_WIRE_69);


b2v_inst39 : static_1
PORT MAP(		 o => SYNTHESIZED_WIRE_57);


b2v_inst4 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_62,
		 b => SYNTHESIZED_WIRE_63,
		 c => SYNTHESIZED_WIRE_22);


b2v_inst40 : static_0
PORT MAP(		 o => SYNTHESIZED_WIRE_59);


b2v_inst5 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_64,
		 b => SYNTHESIZED_WIRE_65,
		 c => SYNTHESIZED_WIRE_10);


b2v_inst6 : gf_sum
PORT MAP(a => SYNTHESIZED_WIRE_77,
		 b => SYNTHESIZED_WIRE_78,
		 c => SYNTHESIZED_WIRE_26);


b2v_inst7 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_69,
		 o => SYNTHESIZED_WIRE_64);


b2v_inst8 : gf_mult
PORT MAP(x => SYNTHESIZED_WIRE_74,
		 y => SYNTHESIZED_WIRE_71,
		 o => SYNTHESIZED_WIRE_54);



END bdf_type;