
library ieee;
use ieee.std_logic_1164.all;

entity manchester_decoder is

	port
	(
		clk		 : in	std_logic;
		data_in	 : in	std_logic;
		reset	 : in	std_logic;
		data_out : out	std_logic;
		s : out std_logic_vector(3 downto 0)
	);
	
end entity;

architecture rtl of manchester_decoder is

	-- Build an enumerated type for the state machine
	type state_type is (s0, s1, s2, s3, s4);
	
	-- Register to hold the current state
	signal state : state_type;

begin
	process (clk, reset)
	begin
		if reset = '1' then
			state <= s0;
		elsif (rising_edge(clk)) then
			-- Determine the next state synchronously, based on
			-- the current state and the input
			case state is
				when s0=>
					if data_in = '1' then
						state <= s2;
					else
						state <= s1;
					end if;
				when s1=>
					if data_in = '1' then
						state <= s3;
					else
						state <= s0;
					end if;
				when s2=>
					if data_in = '1' then
						state <= s0;
					else
						state <= s4;
					end if;
				when s3=>
					if data_in = '1' then
						state <= s2;
					else
						state <= s1;
					end if;
				when s4=>
					if data_in = '1' then
						state <= s2;
					else
						state <= s1;
					end if;
			end case;
			
		end if;
	end process;
	
	process (state)
	begin
		case state is
			when s0=>
				if data_in = '1' then
					data_out <= '1';
					s <= "0000";
				else
					data_out <= '0';
					s <= "0001";
				end if;
			when s1=>
					data_out <= '0';
					s <= "0010";
			when s2=>
					data_out <= '1';
					s <= "0011";
			when s3=>

					s <= "0100";
					data_out <= '0';

			when s4=>
					data_out <= '1';
					s <= "0101";
		end case;
	end process;
	
end rtl;
