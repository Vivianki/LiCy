LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY xor5x1 IS 
	PORT
	(
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		C1 :  IN  STD_LOGIC;
		D1 :  IN  STD_LOGIC;
		E1 :  IN  STD_LOGIC;
		F :  OUT  STD_LOGIC
	);
END xor5x1;

ARCHITECTURE bdf_type OF xor5x1 IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_1 <= A1 XOR B1;


SYNTHESIZED_WIRE_0 <= C1 XOR D1;


SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_0 XOR E1;


F <= SYNTHESIZED_WIRE_1 XOR SYNTHESIZED_WIRE_2;


END bdf_type;